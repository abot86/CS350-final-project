`timescale 1ns / 1ps

module timing_tb;

    Wrapper_tb cpu();
endmodule