module adc_interface();

endmodule